library verilog;
use verilog.vl_types.all;
entity REG4BIT_vlg_vec_tst is
end REG4BIT_vlg_vec_tst;
